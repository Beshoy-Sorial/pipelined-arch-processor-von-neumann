LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
ENTITY reg_file IS
  port(
    clk:in std_logic;
    write_enable:in std_logic;
    read_reg_address_1:in std_logic_vector(2 downto 0);
        read_reg_address_2:in std_logic_vector(2 downto 0);
        write_reg_address:in std_logic_vector(2 downto 0);
        write_data :in std_logic_vector(31 downto 0);
        read_data_1 :out std_logic_vector(31 downto 0);
        read_data_2 :out std_logic_vector(31 downto 0)
        );
end reg_file;

architecture arch_reg_file of reg_file is 
  type type_array is array (0 to 7) of std_logic_vector (31 downto 0);
  signal register_file : type_array:= (others=>(others=>'0'));
begin
  write_process:process(clk)
  begin 
    if rising_edge(clk)then 
      if write_enable = '1' then 
        register_file(to_integer(unsigned(write_reg_address)))<=write_data;
      end if;
    end if ;
  end process;
  
  
  read_process:process(clk)
  begin 
    if falling_edge(clk)then
      read_data_1<= register_file(to_integer(unsigned(read_reg_address_1)));
      read_data_2<=register_file(to_integer(unsigned(read_reg_address_2)));
    end if ;
  end process;

end arch_reg_file;
